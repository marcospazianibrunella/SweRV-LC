// SPDX-License-Identifier: Apache-2.0
// Copyright 2019 Western Digital Corporation or its affiliates.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// all flops call the rvdff flop

/* Understand if I'm in Sim or not */

// synthesis translate_off
`define IN_SIM
// synthesis translate_on

`ifndef IN_SIM
`ifndef VERILATOR
`include "global.svh"
`endif
`endif

module rvdff #( parameter WIDTH=1 )
   (
     input logic [WIDTH-1:0] din,
     input logic           clk,
     input logic                   rst_l,

     output logic [WIDTH-1:0] dout
     );

`ifdef CLOCKGATE
   always @(posedge tb_top.clk) begin
      #0 $strobe("CG: %0t %m din %x dout %x clk %b width %d",$time,din,dout,clk,WIDTH);
   end
`endif

   always_ff @(posedge clk) begin
      if (rst_l == 0)
        dout[WIDTH-1:0] <= 0;
      else
        dout[WIDTH-1:0] <= din[WIDTH-1:0];
   end


endmodule

// rvdff with 2:1 input mux to flop din iff sel==1
module rvdffs #( parameter WIDTH=1 )
   (
     input logic [WIDTH-1:0] din,
     input logic             en,
     input logic           clk,
     input logic                   rst_l,
     output logic [WIDTH-1:0] dout
     );

   rvdff #(WIDTH) dffs (.din((en) ? din[WIDTH-1:0] : dout[WIDTH-1:0]), .*);

endmodule

// rvdff with en and clear
module rvdffsc #( parameter WIDTH=1 )
   (
     input logic [WIDTH-1:0] din,
     input logic             en,
     input logic             clear,
     input logic           clk,
     input logic                   rst_l,
     output logic [WIDTH-1:0] dout
     );

   logic [WIDTH-1:0]          din_new;
   assign din_new = {WIDTH{~clear}} & (en ? din[WIDTH-1:0] : dout[WIDTH-1:0]);
   rvdff #(WIDTH) dffsc (.din(din_new[WIDTH-1:0]), .*);

endmodule

// versions with clock enables .clken to assist in RV_FPGA_OPTIMIZE
module rvdff_fpga #( parameter WIDTH=1 )
   (
     input logic [WIDTH-1:0] din,
     input logic           clk,
     input logic           clken,
     input logic           rawclk,
     input logic           rst_l,
     input logic           scan_mode,

     output logic [WIDTH-1:0] dout
     );

`ifdef RV_FPGA_OPTIMIZE
    rvdffs #(WIDTH) dffs (.clk(rawclk), .en(clken), .*);
`else
    rvdff #(WIDTH)  dff (.*);
`endif



endmodule

// rvdff with 2:1 input mux to flop din iff sel==1
module rvdffs_fpga #( parameter WIDTH=1 )
   (
     input logic [WIDTH-1:0] din,
     input logic             en,
     input logic           clk,
     input logic           clken,
     input logic           rawclk,
     input logic           rst_l,
     input logic           scan_mode,
     output logic [WIDTH-1:0] dout
     );

`ifdef RV_FPGA_OPTIMIZE
   rvdffs #(WIDTH)   dffs (.clk(rawclk), .en(clken & en), .*);
`else
   rvdffs #(WIDTH)   dffs (.*);
`endif

endmodule

// rvdff with en and clear
module rvdffsc_fpga #( parameter WIDTH=1 )
   (
     input logic [WIDTH-1:0] din,
     input logic             en,
     input logic             clear,
     input logic             clk,
     input logic             clken,
     input logic             rawclk,
     input logic             rst_l,
     input logic             scan_mode,
     output logic [WIDTH-1:0] dout
     );

`ifdef RV_FPGA_OPTIMIZE
   rvdffs  #(WIDTH)   dffs  (.clk(rawclk), .din(din[WIDTH-1:0] & {WIDTH{~clear}}),.en((en | clear) & clken), .*);
`else
   rvdffsc #(WIDTH)   dffsc (.*);
`endif

endmodule


module `TEC_RV_ICG
  (
   input logic TE, E, CP,
   output Q
   );

   logic  en_ff;
   logic  enable;

   assign      enable = E | TE;

`ifdef VERILATOR
   always @(negedge CP) begin
      en_ff <= enable;
   end
`else
   always @(CP, enable) begin
      if(!CP)
        en_ff = enable;
   end
`endif
   assign Q = CP & en_ff;

endmodule

`ifndef RV_FPGA_OPTIMIZE
module rvclkhdr
  (
   input  logic en,
   input  logic clk,
   input  logic scan_mode,
   output logic l1clk
   );

   logic        TE;
   assign       TE = scan_mode;

   `TEC_RV_ICG clkhdr ( .*, .E(en), .CP(clk), .Q(l1clk));

endmodule // rvclkhdr
`endif

module rvoclkhdr
  (
   input  logic en,
   input  logic clk,
   input  logic scan_mode,
   output logic l1clk
   );

   logic        TE;
   assign       TE = scan_mode;

`ifdef RV_FPGA_OPTIMIZE
   assign l1clk = clk;
`else
   `TEC_RV_ICG rvclkhdr ( .*, .E(en), .CP(clk), .Q(l1clk));
`endif

endmodule

module rvdffe #( parameter WIDTH=1, parameter OVERRIDE=0 )
   (
     input  logic [WIDTH-1:0] din,
     input  logic           en,
     input  logic           clk,
     input  logic           rst_l,
     input  logic             scan_mode,
     output logic [WIDTH-1:0] dout
     );

   logic                      l1clk;


`ifndef PHYSICAL
   if (WIDTH >= 8 || OVERRIDE==1) begin: genblock
`endif

`ifdef RV_FPGA_OPTIMIZE
      rvdffs #(WIDTH) dff ( .* );
`else
      rvclkhdr clkhdr ( .* );
      rvdff #(WIDTH) dff (.*, .clk(l1clk));
`endif

`ifndef PHYSICAL
   end
   else
      $error("%m: rvdffe width must be >= 8");
`endif


endmodule // rvdffe

module rvsyncss #(parameter WIDTH = 251)
   (
     input  logic                 clk,
     input  logic                 rst_l,
     input  logic [WIDTH-1:0]     din,
     output logic [WIDTH-1:0]     dout
     );

   logic [WIDTH-1:0]              din_ff1;

   rvdff #(WIDTH) sync_ff1  (.*, .din (din[WIDTH-1:0]),     .dout(din_ff1[WIDTH-1:0]));
   rvdff #(WIDTH) sync_ff2  (.*, .din (din_ff1[WIDTH-1:0]), .dout(dout[WIDTH-1:0]));

endmodule // rvsyncss

module rvlsadder #(parameter XLEN = 64)
  (
    input logic [XLEN-1:0] rs1,
    input logic [11:0] offset,

    output logic [XLEN-1:0] dout
    );

   logic                cout;
   logic                sign;

   logic [XLEN-1:12]        rs1_inc;
   logic [XLEN-1:12]        rs1_dec;

   assign {cout,dout[11:0]} = {1'b0,rs1[11:0]} + {1'b0,offset[11:0]};

   assign rs1_inc[XLEN-1:12] = rs1[XLEN-1:12] + 1;

   assign rs1_dec[XLEN-1:12] = rs1[XLEN-1:12] - 1;

   assign sign = offset[11];

   assign dout[XLEN-1:12] = ({XLEN-12{  sign ^~  cout}} &     rs1[XLEN-1:12]) |
                        ({XLEN-12{ ~sign &   cout}}  & rs1_inc[XLEN-1:12]) |
                        ({XLEN-12{  sign &  ~cout}}  & rs1_dec[XLEN-1:12]);

endmodule // rvlsadder

// assume we only maintain pc[31:1] in the pipe

module rvbradder
  (
    input [31:1] pc,
    input [12:1] offset,

    output [31:1] dout
    );

   logic          cout;
   logic          sign;

   logic [31:13]  pc_inc;
   logic [31:13]  pc_dec;

   assign {cout,dout[12:1]} = {1'b0,pc[12:1]} + {1'b0,offset[12:1]};

   assign pc_inc[31:13] = pc[31:13] + 1;

   assign pc_dec[31:13] = pc[31:13] - 1;

   assign sign = offset[12];


   assign dout[31:13] = ({19{  sign ^~  cout}} &     pc[31:13]) |
                        ({19{ ~sign &   cout}}  & pc_inc[31:13]) |
                        ({19{  sign &  ~cout}}  & pc_dec[31:13]);


endmodule // rvbradder


// 2s complement circuit
module rvtwoscomp #( parameter WIDTH=32 )
   (
     input logic [WIDTH-1:0] din,

     output logic [WIDTH-1:0] dout
     );

   logic [WIDTH-1:1]          dout_temp;   // holding for all other bits except for the lsb. LSB is always din

   genvar                     i;

   for ( i = 1; i < WIDTH; i++ )  begin : flip_after_first_one
      assign dout_temp[i] = (|din[i-1:0]) ? ~din[i] : din[i];
   end : flip_after_first_one

   assign dout[WIDTH-1:0]  = { dout_temp[WIDTH-1:1], din[0] };

endmodule  // 2'scomp

// find first
module rvfindfirst1 #( parameter WIDTH=32, SHIFT=$clog2(WIDTH) )
   (
     input logic [WIDTH-1:0] din,

     output logic [SHIFT-1:0] dout
     );
   logic                      done;

   always_comb begin
      dout[SHIFT-1:0] = {SHIFT{1'b0}};
      done    = 1'b0;

      for ( int i = WIDTH-1; i > 0; i-- )  begin : find_first_one
         done |= din[i];
         dout[SHIFT-1:0] += done ? 1'b0 : 1'b1;
      end : find_first_one
   end
endmodule // rvfindfirst1

module rvfindfirst1hot #( parameter WIDTH=32 )
   (
     input logic [WIDTH-1:0] din,

     output logic [WIDTH-1:0] dout
     );
   logic                      done;

   always_comb begin
      dout[WIDTH-1:0] = {WIDTH{1'b0}};
      done    = 1'b0;
      for ( int i = 0; i < WIDTH; i++ )  begin : find_first_one
         dout[i] = ~done & din[i];
         done   |= din[i];
      end : find_first_one
   end
endmodule // rvfindfirst1hot

// mask and match function matches bits after finding the first 0 position
// find first starting from LSB. Skip that location and match the rest of the bits
module rvmaskandmatch #( parameter WIDTH=32 )
   (
     input  logic [WIDTH-1:0] mask,     // this will have the mask in the lower bit positions
     input  logic [WIDTH-1:0] data,     // this is what needs to be matched on the upper bits with the mask's upper bits
     input  logic             masken,   // when 1 : do mask. 0 : full match
     output logic             match
     );

   logic [WIDTH-1:0]          matchvec;
   logic                      masken_or_fullmask;

   assign masken_or_fullmask = masken &  ~(&mask[WIDTH-1:0]);

   assign matchvec[0]        = masken_or_fullmask | (mask[0] == data[0]);
   genvar                     i;

   for ( i = 1; i < WIDTH; i++ )  begin : match_after_first_zero
      assign matchvec[i] = (&mask[i-1:0] & masken_or_fullmask) ? 1'b1 : (mask[i] == data[i]);
   end : match_after_first_zero

   assign match  = &matchvec[WIDTH-1:0];    // all bits either matched or were masked off

endmodule // rvmaskandmatch

module rvbtb_tag_hash (
                       input logic [31:1] pc,
                       output logic [`RV_BTB_BTAG_SIZE-1:0] hash
                       );
`ifndef RV_BTB_BTAG_FOLD
    assign hash = {(pc[`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE+`RV_BTB_BTAG_SIZE+`RV_BTB_BTAG_SIZE:`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE+`RV_BTB_BTAG_SIZE+1] ^
                   pc[`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE+`RV_BTB_BTAG_SIZE:`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE+1] ^
                   pc[`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE:`RV_BTB_ADDR_HI+1])};
`else
    assign hash = {(
                   pc[`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE+`RV_BTB_BTAG_SIZE:`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE+1] ^
                   pc[`RV_BTB_ADDR_HI+`RV_BTB_BTAG_SIZE:`RV_BTB_ADDR_HI+1])};
`endif

//  assign hash = {pc[`RV_BTB_ADDR_HI+1],(pc[`RV_BTB_ADDR_HI+13:`RV_BTB_ADDR_HI+10] ^
//                                       pc[`RV_BTB_ADDR_HI+9:`RV_BTB_ADDR_HI+6] ^
//                                       pc[`RV_BTB_ADDR_HI+5:`RV_BTB_ADDR_HI+2])};

endmodule

module rvbtb_addr_hash (
                        input logic [31:1] pc,
                        output logic [`RV_BTB_ADDR_HI:`RV_BTB_ADDR_LO] hash
                        );

   assign hash[`RV_BTB_ADDR_HI:`RV_BTB_ADDR_LO] = pc[`RV_BTB_INDEX1_HI:`RV_BTB_INDEX1_LO] ^

`ifndef RV_BTB_FOLD2_INDEX_HASH
                                                  pc[`RV_BTB_INDEX2_HI:`RV_BTB_INDEX2_LO] ^
`endif

                                                  pc[`RV_BTB_INDEX3_HI:`RV_BTB_INDEX3_LO];

endmodule

module rvbtb_ghr_hash (
                       input logic [`RV_BTB_ADDR_HI:`RV_BTB_ADDR_LO] hashin,
                       input logic [`RV_BHT_GHR_RANGE] ghr,
                       output logic [`RV_BHT_ADDR_HI:`RV_BHT_ADDR_LO] hash
                       );

   // The hash function is too complex to write in verilog for all cases.
   // The config script generates the logic string based on the bp config.
   assign hash[`RV_BHT_ADDR_HI:`RV_BHT_ADDR_LO] = `RV_BHT_HASH_STRING;

endmodule


// Check if the S_ADDR <= addr < E_ADDR
module rvrangecheck  #(CCM_SADR = 32'h0,
                       CCM_SIZE  = 128) (
   input  logic [31:0]   addr,                             // Address to be checked for range
   output logic          in_range,                            // S_ADDR <= start_addr < E_ADDR
   output logic          in_region
);

   localparam REGION_BITS = 4;
   localparam MASK_BITS = 10 + $clog2(CCM_SIZE);

   logic [31:0]          start_addr;
   logic [3:0]           region;

   assign start_addr[31:0]        = CCM_SADR;
   assign region[REGION_BITS-1:0] = start_addr[31:(32-REGION_BITS)];

   assign in_region = (addr[31:(32-REGION_BITS)] == region[REGION_BITS-1:0]);
   if (CCM_SIZE  == 48)
    assign in_range  = (addr[31:MASK_BITS] == start_addr[31:MASK_BITS]) & ~(&addr[MASK_BITS-1 : MASK_BITS-2]);
   else
    assign in_range  = (addr[31:MASK_BITS] == start_addr[31:MASK_BITS]);

endmodule  // rvrangechecker

// 16 bit even parity generator
module rveven_paritygen #(WIDTH = 16)  (
                                         input  logic [WIDTH-1:0]  data_in,         // Data
                                         output logic              parity_out       // generated even parity
                                         );

   assign  parity_out =  ^(data_in[WIDTH-1:0]) ;

endmodule  // rveven_paritygen

module rveven_paritycheck #(WIDTH = 16)  (
                                           input  logic [WIDTH-1:0]  data_in,         // Data
                                           input  logic              parity_in,
                                           output logic              parity_err       // Parity error
                                           );

   assign  parity_err =  ^(data_in[WIDTH-1:0]) ^ parity_in ;

endmodule  // rveven_paritycheck

module rvecc_encode  (
                      input [63:0] din,
                      output [7:0] ecc_out
                      );
logic [5:0] ecc_out_temp;

   assign ecc_out_temp[0] = din[0]^din[1]^din[3]^din[4]^din[6]^din[8]^din[10]^din[11]^din[13]^din[15]^din[17]^din[19]^din[21]^din[23]^din[25]^din[26]^din[28]^din[30]
                            ^din[32]^din[34]^din[36]^din[38]^din[40]^din[42]^din[44]^din[46]^din[48]^din[50]^din[52]^din[54]^din[56]^din[57]^din[59]^din[61]^din[63];

   assign ecc_out_temp[1] = din[0]^din[2]^din[3]^din[5]^din[6]^din[9]^din[10]^din[12]^din[13]^din[16]^din[17]^din[20]^din[21]^din[24]^din[25]^din[27]^din[28]^din[31]
                            ^din[32]^din[32]^din[36]^din[39]^din[40]^din[43]^din[44]^din[47]^din[48]^din[51]^din[52]^din[55]^din[56]^din[58]^din[59]^din[62]^din[63];

   assign ecc_out_temp[2] = din[1]^din[2]^din[3]^din[7]^din[8]^din[9]^din[10]^din[14]^din[15]^din[16]^din[17]^din[22]^din[23]^din[24]^din[25]^din[29]^din[30]^din[31]
                            ^din[32]^din[37]^din[38]^din[39]^din[40]^din[45]^din[46]^din[47]^din[48]^din[53]^din[54]^din[55]^din[56]^din[60]^din[61]^din[62]^din[63];

   assign ecc_out_temp[3] = din[4]^din[5]^din[6]^din[7]^din[8]^din[9]^din[10]^din[18]^din[19]^din[20]^din[21]^din[22]^din[23]^din[24]^din[25]
                            ^din[33]^din[34]^din[35]^din[36]^din[37]^din[38]^din[39]^din[40]^din[49]^din[50]^din[51]^din[52]^din[53]^din[54]^din[55]^din[56];

   assign ecc_out_temp[4] = din[11]^din[12]^din[13]^din[14]^din[15]^din[16]^din[17]^din[18]^din[19]^din[20]^din[21]^din[22]^din[23]^din[24]^din[25]
                            ^din[41]^din[42]^din[43]^din[44]^din[45]^din[46]^din[47]^din[48]^din[49]^din[50]^din[51]^din[52]^din[53]^din[54]^din[55]^din[56];

   assign ecc_out_temp[5] = ^din[56:26];
   
   assign ecc_out_temp[6] = ^din[63:57];

   assign ecc_out[7:0] = {(^din[63:0])^(^ecc_out_temp[6:0]),ecc_out_temp[6:0]};

endmodule // rvecc_encode

module rvecc_decode  (
                      input         en,
                      input [63:0]  din,
                      input [7:0]   ecc_in,
                      input         sed_ded,    // only do detection and no correction. Used for the I$
                      output [63:0] dout,
                      output [7:0]  ecc_out,
                      output        single_ecc_error,
                      output        double_ecc_error

                      );

   logic [7:0]                      ecc_check;
   logic [63:0]                     error_mask;
   logic [71:0]                     din_plus_parity, dout_plus_parity;

   // Syndrome Generation
   assign ecc_check[0] = ecc_in[0]^din[0]^din[1]^din[3]^din[4]^din[6]^din[8]^din[10]^din[11]^din[13]^din[15]^din[17]^din[19]^din[21]^din[23]^din[25]^din[26]^din[28]^din[30]
   ^din[32]^din[34]^din[36]^din[38]^din[40]^din[42]^din[44]^din[46]^din[48]^din[50]^din[52]^din[54]^din[56]^din[57]^din[59]^din[61]^din[63];

   assign ecc_check[1] = ecc_in[1]^din[0]^din[2]^din[3]^din[5]^din[6]^din[9]^din[10]^din[12]^din[13]^din[16]^din[17]^din[20]^din[21]^din[24]^din[25]^din[27]^din[28]^din[31]
   ^din[32]^din[32]^din[36]^din[39]^din[40]^din[43]^din[44]^din[47]^din[48]^din[51]^din[52]^din[55]^din[56]^din[58]^din[59]^din[62]^din[63];

   assign ecc_check[2] = ecc_in[2]^din[1]^din[2]^din[3]^din[7]^din[8]^din[9]^din[10]^din[14]^din[15]^din[16]^din[17]^din[22]^din[23]^din[24]^din[25]^din[29]^din[30]^din[31]
   ^din[32]^din[37]^din[38]^din[39]^din[40]^din[45]^din[46]^din[47]^din[48]^din[53]^din[54]^din[55]^din[56]^din[60]^din[61]^din[62]^din[63];

   assign ecc_check[3] = ecc_in[3]^din[4]^din[5]^din[6]^din[7]^din[8]^din[9]^din[10]^din[18]^din[19]^din[20]^din[21]^din[22]^din[23]^din[24]^din[25]
   ^din[33]^din[34]^din[35]^din[36]^din[37]^din[38]^din[39]^din[40]^din[49]^din[50]^din[51]^din[52]^din[53]^din[54]^din[55]^din[56];

   assign ecc_check[4] = ecc_in[4]^din[11]^din[12]^din[13]^din[14]^din[15]^din[16]^din[17]^din[18]^din[19]^din[20]^din[21]^din[22]^din[23]^din[24]^din[25]
   ^din[41]^din[42]^din[43]^din[44]^din[45]^din[46]^din[47]^din[48]^din[49]^din[50]^din[51]^din[52]^din[53]^din[54]^din[55]^din[56];

   assign ecc_check[5] = ecc_in[5]^(^din[56:26]);
   
   assign ecc_check[6] = ecc_in[6]^(^din[63:57]);

   // This is the parity bit
   assign ecc_check[7] = ((^din[63:0])^(^ecc_in[6:0])) & ~sed_ded;

   assign single_ecc_error = en & (ecc_check[7:0] != 0) & ecc_check[7];   // this will never be on for sed_ded
   assign double_ecc_error = en & (ecc_check[7:0] != 0) & ~ecc_check[7];  // all errors in the sed_ded case will be recorded as DE

   //// Generate the mask for error correctiong
   always @(*)begin 
         case (ecc_check)
            8'b10000011 :
                     begin
                        error_mask <= 64'h0000000000000001 ; // 0
                     end
            8'b10000101 :
                     begin
                        error_mask <= 64'h0000000000000002 ; // 1			
                     end
            8'b10000110 :
                     begin
                        error_mask <= 64'h0000000000000004 ; // 2			
                     end
            8'b10000111 :
                     begin
                        error_mask <= 64'h0000000000000008 ; // 3
                     end
            8'b10001001 :
                     begin
                        error_mask <= 64'h0000000000000010 ; // 4
                     end
            8'b10001010 :
                     begin
                        error_mask <= 64'h0000000000000020 ; // 5
                     end
            8'b10001011 :
                     begin
                        error_mask <= 64'h0000000000000040 ; // 6
                     end
            8'b10001100 :
                     begin
                        error_mask <= 64'h0000000000000080 ; // 7
                     end
            8'b10001101 :
                     begin
                        error_mask <= 64'h0000000000000100 ; // 8
                     end
            8'b10001110 :
                     begin
                        error_mask <= 64'h0000000000000200 ; // 9
                     end
            8'b10001111 :
                     begin
                        error_mask <= 64'h0000000000000400 ; // 10
                     end
            8'b10010001 :
                     begin
                        error_mask <= 64'h0000000000000800 ; // 11
                     end
            8'b10010010 :
                     begin
                        error_mask <= 64'h0000000000001000 ; // 12
                     end
            8'b10010011 :
                     begin
                        error_mask <= 64'h0000000000002000 ; // 13
                     end
            8'b10010100 :
                     begin
                        error_mask <= 64'h0000000000004000 ; // 14
                     end
            8'b10010101 :
                     begin
                        error_mask <= 64'h0000000000008000 ; // 15
                     end
            8'b10010110 :
                     begin
                        error_mask <= 64'h0000000000010000 ; // 16
                     end
            8'b10010111 :
                     begin
                        error_mask <= 64'h0000000000020000 ; // 17
                     end
            8'b10011000 :
                     begin
                        error_mask <= 64'h0000000000040000 ; // 18
                     end
            8'b10011001 :
                     begin
                        error_mask <= 64'h0000000000080000 ; // 19
                     end
            8'b10011010 :
                     begin
                        error_mask <= 64'h0000000000100000 ; // 20
                     end
            8'b10011011 :
                     begin
                        error_mask <= 64'h0000000000200000 ; // 21
                     end
            8'b10011100 :
                     begin
                        error_mask <= 64'h0000000000400000 ; // 22
                     end
            8'b10011101 :
                     begin
                        error_mask <= 64'h0000000000800000 ; // 23
                     end
            8'b10011110 :
                     begin
                        error_mask <= 64'h0000000001000000 ; // 24
                     end
            8'b10011111 :
                     begin
                        error_mask <= 64'h0000000002000000 ; // 25
                     end
            8'b10100001 :
                     begin
                        error_mask <= 64'h0000000004000000 ; // 26
                     end
            8'b10100010 :
                     begin
                        error_mask <= 64'h0000000008000000 ; // 27
                     end
            8'b10100011 :
                     begin
                        error_mask <= 64'h0000000010000000 ; // 28
                     end
            8'b10100100 :
                     begin
                        error_mask <= 64'h0000000020000000 ; // 29
                     end
            8'b10100101 :
                     begin
                        error_mask <= 64'h0000000040000000 ; // 30
                     end
            8'b10100110 :
                     begin
                        error_mask <= 64'h0000000080000000 ; // 31
                     end
            8'b10100111 :
                     begin
                        error_mask <= 64'h0000000100000000 ; // 32
                     end
            8'b10101000 :
                     begin
                        error_mask <= 64'h0000000200000000 ; // 33
                     end
            8'b10101001 :
                     begin
                        error_mask <= 64'h0000000400000000 ; // 34
                     end
            8'b10101010 :
                     begin
                        error_mask <= 64'h0000000800000000 ; // 35
                     end
            8'b10101011 :
                     begin
                        error_mask <= 64'h0000001000000000 ; // 36
                     end
            8'b10101100 :
                     begin
                        error_mask <= 64'h0000002000000000 ; // 37
                     end
            8'b10101101 :
                     begin
                        error_mask <= 64'h0000004000000000 ; // 38
                     end
            8'b10101110 :
                     begin
                        error_mask <= 64'h0000008000000000 ; // 39
                     end
            8'b10101111 :
                     begin
                        error_mask <= 64'h0000010000000000 ; // 40
                     end
            8'b10110000 :
                     begin
                        error_mask <= 64'h0000020000000000 ; // 41
                     end
            8'b10110001 :
                     begin
                        error_mask <= 64'h0000040000000000 ; // 42
                     end
            8'b10110010 :
                     begin
                        error_mask <= 64'h0000080000000000 ; // 43
                     end
            8'b10110011 :
                     begin
                        error_mask <= 64'h0000100000000000 ; // 44
                     end
            8'b10110100 :
                     begin
                        error_mask <= 64'h0000200000000000 ; // 45
                     end
            8'b10110101 :
                     begin
                        error_mask <= 64'h0000400000000000 ; // 46
                     end
            8'b10110110 :
                     begin
                        error_mask <= 64'h0000800000000000 ; // 47
                     end
            8'b10110111 :
                     begin
                        error_mask <= 64'h0001000000000000 ; // 48
                     end
            8'b10111000 :
                     begin
                        error_mask <= 64'h0002000000000000 ; // 49
                     end
            8'b10111001 :
                     begin
                        error_mask <= 64'h0004000000000000 ; // 50
                     end
            8'b10111010 :
                     begin
                        error_mask <= 64'h0008000000000000 ; // 51
                     end
            8'b10111011 :
                     begin
                        error_mask <= 64'h0010000000000000 ; // 52
                     end
            8'b10111100 :
                     begin
                        error_mask <= 64'h0020000000000000 ; // 53
                     end
            8'b10111101 :
                     begin
                        error_mask <= 64'h0040000000000000 ; // 54
                     end
            8'b10111110 :
                     begin
                        error_mask <= 64'h0080000000000000 ; // 55
                     end
            8'b10111111 :
                     begin
                        error_mask <= 64'h0100000000000000 ; // 56
                     end
            8'b11000001 :
                     begin
                        error_mask <= 64'h0200000000000000 ; // 57
                     end
            8'b11000010 :
                     begin
                        error_mask <= 64'h0400000000000000 ; // 58
                     end
            8'b11000011 :
                     begin
                        error_mask <= 64'h0800000000000000 ; // 59
                     end
            8'b11000100 :
                     begin
                        error_mask <= 64'h1000000000000000 ; // 60
                     end
            8'b11000101 :
                     begin
                        error_mask <= 64'h2000000000000000 ; // 61
                     end
            8'b11000110 :
                     begin
                        error_mask <= 64'h4000000000000000 ; // 62
                     end
            8'b11000111 :
                     begin
                        error_mask <= 64'h8000000000000000 ; // 63	
                     end
            default :
                     begin
                        error_mask <= 64'h0000000000000000 ; 
                     end
         endcase 
   end 

   // Generate the corrected data
   assign dout[63:0]             = mask ^ din;
   assign ecc_out[7:0]           = {(dout_plus_parity[38] ^ (ecc_check[7:0] == 8'b1000_0000)), dout_plus_parity[31], dout_plus_parity[15], dout_plus_parity[7], dout_plus_parity[3], dout_plus_parity[1:0]};

endmodule // rvecc_decode
